LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY uc IS
PORT	(	F		:	IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			EnA, EnB, InvA, InvB, C0, O1, O0		:	OUT STD_LOGIC);
END uc;
ARCHITECTURE funcionamento OF uc IS

SIGNAL D	:	STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
	WITH F SELECT
		D <=  "00000001" WHEN "000",
				"00000010" WHEN "001",   	
				"00000100" WHEN "010", 
				"00001000" WHEN "011",
				"00010000" WHEN "100",
				"00100000" WHEN "101",
				"01000000" WHEN "110",
				"10000000" WHEN "111",
				"00000000" WHEN OTHERS;
	EnA <= D(1) OR D(2) OR D(3);
	EnB <= D(1) OR D(2) OR D(3);
	InvB <= D(1) OR D(7);
	InvA <= D(2);
	C0 <= D(1) OR D(2);
	O0 <= D(4) OR D(5);
	O1 <= D(4) OR D(6);
	
	
END funcionamento;