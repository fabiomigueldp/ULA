LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FA IS
PORT	(	Ai, Bi, Cin		:	IN STD_LOGIC;
			Cout, Si			:	OUT STD_LOGIC);
END FA;

ARCHITECTURE sumbit OF FA IS
SIGNAL X:	STD_LOGIC;
BEGIN
	X <= Ai XOR Bi;
	Si <= X XOR Cin;
	Cout <= (Ai AND Bi) OR (X AND Cin);
END sumbit;