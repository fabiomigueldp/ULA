LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX IS
PORT ( Re,Rxor,Rou,Rs: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O1, O0 : IN STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END MUX;

ARCHITECTURE multi OF MUX IS
SIGNAL O : STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN 
	O <= O1 & O0;
	WITH  O SELECT
	S <= Rs WHEN "00",
		  Rou WHEN "01",
		  Re WHEN "10",
		  Rxor WHEN "11";
END multi;