LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ULA IS
PORT   (
		A,B : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		F : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		sS, dSd, dSu: OUT STD_LOGIC_VECTOR(0 TO 6);
		E : OUT STD_LOGIC);
END ULA;

ARCHITECTURE arquitetura OF ULA IS
	SIGNAL EnA, EnB, InvA, InvB, C0 : STD_LOGIC;
	SIGNAL Re, Rxor, Rou, Rs : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL O1, O0 : STD_LOGIC;
	SIGNAL S : STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	COMPONENT ul
	PORT	(	A,B		:	IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			Re, Rxor, Rou		:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT MUX
	PORT ( Re,Rxor,Rou,Rs: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O1, O0 : IN STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT somasub
	PORT	(	A,B		:	IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				EnA, EnB, InvA, InvB, C0	:	IN STD_LOGIC;
				E		:	OUT STD_LOGIC;
				Rs		:  OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT uc
	PORT	(	F		:	IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			EnA, EnB, InvA, InvB, C0, O1, O0		:	OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT DISPLAY
	PORT (valor			: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			sinal			: IN STD_LOGIC;
			digS, dig1, dig0	: OUT STD_LOGIC_VECTOR(0 TO 6));	
	END COMPONENT;
	
BEGIN 

	UC0 : uc PORT MAP (F, EnA, EnB, InvA, InvB, C0, O1, O0);
	UA0 : somasub PORT MAP (A, B, EnA, EnB, InvA, InvB, C0, E, Rs);
	UL0 : ul PORT MAP (A,B, Re, Rxor, Rou);
	MUX0 : MUX PORT MAP (Re, Rxor, Rou, Rs, O1, O0, S);
	DSPS : DISPLAY PORT MAP (S, '1', sS, dSd, dSu);

END arquitetura;