LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ULA IS
PORT   (
		A,B : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		F : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		E : OUT STD_LOGIC);
END ULA;

ARCHITECTURE arquitetura OF ULA IS
	SIGNAL EnA, EnB, InvA, InvB, C0 : STD_LOGIC;
	SIGNAL Re, Rxor, Rou, Rs : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL O1, O0 : STD_LOGIC;
	SIGNAL S : STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	COMPONENT MUX
	PORT ( Re,Rxor,Rou,Rs: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O1, O0 : IN STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT somasub
	PORT	(	A,B		:	IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				EnA, EnB, InvA, InvB, C0	:	IN STD_LOGIC;
				E		:	OUT STD_LOGIC;
				Rs		:  OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT uc
	PORT	(	F		:	IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			EnA, EnB, InvA, InvB, C0, O1, O0		:	OUT STD_LOGIC);
	END COMPONENT;
	
BEGIN 
	Re <= (OTHERS => 'X');
	Rxor <= (OTHERS => 'X');
	Rou <= (OTHERS => 'X');

	UC0 : uc PORT MAP (F, EnA, EnB, InvA, InvB, C0, O1, O0);
	UA0 : somasub PORT MAP (A, B, EnA, EnB, InvA, InvB, C0, E, Rs);
	MUX0 : MUX PORT MAP (Re, Rxor, Rou, Rs, O1, O0, S);

END arquitetura;